`timescale 1ns / 1ps

module i2c_bit_controller_tb;
	
endmodule
