`timescale 1ns/1ps

module i2c_master_controller (
	
);

endmodule

